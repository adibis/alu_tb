`ifndef ALU_TEST_PKG__SV
`define ALU_TEST_PKG__SV

package alu_test_pkg;

    import uvm_pkg::*;
    import alu_pkg::*;
    import env_pkg::*;


    `include "uvm_macros.svh"

    `include "alu_base_test.sv"

endpackage: alu_test_pkg
`endif
