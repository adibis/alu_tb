`ifndef ALU_SEQ_LIST__SV
`define ALU_SEQ_LIST__SV

import uvm_pkg::*;

`include "uvm_macros.svh"

`include "alu_base_seq.sv"

`endif
