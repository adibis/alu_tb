`ifndef ALU_PKG__SV
`define ALU_PKG__SV

package alu_pkg;

    import uvm_pkg::*;

    `include "uvm_macros.svh"

    `include "alu_base_seq_item.sv"
    `include "alu_driver.sv"
    `include "alu_monitor.sv"
    `include "alu_agent.sv"

    `include "alu_seq_list.sv"

endpackage: alu_pkg
`endif
